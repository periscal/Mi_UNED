-- ================================
library IEEE;
use IEEE.std_logic_1164.all;

entity fun2 is
    port(   F28,F29,F30,F31 : out  std_logic;
            A,B,C,D,E       : in   std_logic);
end entity fun2;