-- ================================
-- entity del circuito
-- fichero: fun1.vhd
library IEEE;
use IEEE.std_logic_1164.all;

entity fun1 is port
	(F,G	: out std_logic;
	 A,B,C	: in  std_logic);
end entity fun1;
--=================================